import "DPI-C" function int ebreak();
module EbreakBox ();
ebreak();
endmodule
    
