
import "DPI-C" function void set_gpr_ptr(input logic [63:0] a []);
module Difftest (difftest_gpr_0,difftest_gpr_1,difftest_gpr_2,difftest_gpr_3,difftest_gpr_4,difftest_gpr_5,difftest_gpr_6,difftest_gpr_7,difftest_gpr_8,difftest_gpr_9,difftest_gpr_10,difftest_gpr_11,difftest_gpr_12,difftest_gpr_13,difftest_gpr_14,difftest_gpr_15,difftest_gpr_16,difftest_gpr_17,difftest_gpr_18,difftest_gpr_19,difftest_gpr_20,difftest_gpr_21,difftest_gpr_22,difftest_gpr_23,difftest_gpr_24,difftest_gpr_25,difftest_gpr_26,difftest_gpr_27,difftest_gpr_28,difftest_gpr_29,difftest_gpr_30,difftest_gpr_31,difftest_gpr_32);
 input [63:0] difftest_gpr_0;
 input [63:0] difftest_gpr_1;
 input [63:0] difftest_gpr_2;
 input [63:0] difftest_gpr_3;
 input [63:0] difftest_gpr_4;
 input [63:0] difftest_gpr_5;
 input [63:0] difftest_gpr_6;
 input [63:0] difftest_gpr_7;
 input [63:0] difftest_gpr_8;
 input [63:0] difftest_gpr_9;
 input [63:0] difftest_gpr_10;
 input [63:0] difftest_gpr_11;
 input [63:0] difftest_gpr_12;
 input [63:0] difftest_gpr_13;
 input [63:0] difftest_gpr_14;
 input [63:0] difftest_gpr_15;
 input [63:0] difftest_gpr_16;
 input [63:0] difftest_gpr_17;
 input [63:0] difftest_gpr_18;
 input [63:0] difftest_gpr_19;
 input [63:0] difftest_gpr_20;
 input [63:0] difftest_gpr_21;
 input [63:0] difftest_gpr_22;
 input [63:0] difftest_gpr_23;
 input [63:0] difftest_gpr_24;
 input [63:0] difftest_gpr_25;
 input [63:0] difftest_gpr_26;
 input [63:0] difftest_gpr_27;
 input [63:0] difftest_gpr_28;
 input [63:0] difftest_gpr_29;
 input [63:0] difftest_gpr_30;
 input [63:0] difftest_gpr_31;
 input [63:0] difftest_gpr_32;
 Wire [63:0] rf[32:0];
 assign rf[0]=difftest_gpr_0;
 assign rf[1]=difftest_gpr_1;
 assign rf[2]=difftest_gpr_2;
 assign rf[3]=difftest_gpr_3;
 assign rf[4]=difftest_gpr_4;
 assign rf[5]=difftest_gpr_5;
 assign rf[6]=difftest_gpr_6;
 assign rf[7]=difftest_gpr_7;
 assign rf[8]=difftest_gpr_8;
 assign rf[9]=difftest_gpr_9;
 assign rf[10]=difftest_gpr_10;
 assign rf[11]=difftest_gpr_11;
 assign rf[12]=difftest_gpr_12;
 assign rf[13]=difftest_gpr_13;
 assign rf[14]=difftest_gpr_14;
 assign rf[15]=difftest_gpr_15;
 assign rf[16]=difftest_gpr_16;
 assign rf[17]=difftest_gpr_17;
 assign rf[18]=difftest_gpr_18;
 assign rf[19]=difftest_gpr_19;
 assign rf[20]=difftest_gpr_20;
 assign rf[21]=difftest_gpr_21;
 assign rf[22]=difftest_gpr_22;
 assign rf[23]=difftest_gpr_23;
 assign rf[24]=difftest_gpr_24;
 assign rf[25]=difftest_gpr_25;
 assign rf[26]=difftest_gpr_26;
 assign rf[27]=difftest_gpr_27;
 assign rf[28]=difftest_gpr_28;
 assign rf[29]=difftest_gpr_29;
 assign rf[30]=difftest_gpr_30;
 assign rf[31]=difftest_gpr_31;
 assign rf[32]=difftest_gpr_32;
 initial set_gpr_ptr(rf);
endmodule
    