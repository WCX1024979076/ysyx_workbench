import "DPI-C" function integer \$ebreak;
module EbreakBox ();
$ebreak();
endmodule
    
