import "DPI-C" function void ebreak();
module EbreakBox ();
ebreak();
endmodule
    
