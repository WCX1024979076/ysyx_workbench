
 import "DPI-C" function void ebreak();
 module EbreakBox ();
 function ebreak_fun;
 ebreak();
 end
 endmodule
    